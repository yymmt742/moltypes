netcdf compound_datasize_test2 {
types:
  compound cmpd1 {
    int lat ;
    int lon ;
    int id ;
    uint64 time ;
    int temperature ;
  }; // cmpd1
  compound nested {
    int field1 ;
    int field2 ;
    cmpd1 nested(2) ;
    uint64 field3 ;
    int field4 ;
  }; // nested
dimensions:
	n = UNLIMITED ; // (2 currently)
variables:
	nested scalar ;
	nested array(n) ;
data:

 scalar = 
    {40, -105, {{39, -104, 1111, 7776000, 15}, {39, -104, 1111, 7776000, 15}}, 542932516829005, 17} ;

 array = 
    {40, -105, {{39, -104, 1111, 7776000, 15}, {39, -104, 1111, 7776000, 15}}, 542932516829005, 17}, 
    {40, -105, {{39, -104, 1111, 7776000, 15}, {39, -104, 1111, 7776000, 15}}, 542932516829005, 17} ;
}
