netcdf tst_grp_rename {

types:
  int(*) vlen_t;

dimensions:
  d2 = 2;

variables:
  vlen_t v1(d2);

group: inner {

  types:
    compound c_t { int f1; float f2; };

  dimensions:
    d3 = 3;

  variables:
    c_t vc(d3);

  group: inner_inner {
    dimensions:
      d3 = 4;
  }
}
}
