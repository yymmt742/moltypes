netcdf compound_datasize_test {
types:
  compound obs_t {
    float lat ;
    float lon ;
    string stid ;
    double time ;
    float temperature ;
  }; // obs_t
dimensions:
	n = UNLIMITED ; // (2 currently)
variables:
	obs_t obs(n) ;
data:

 obs = {39.9, -104.9, "KDEN", 7776000, 15}, {40, -105, "KBOU", 7776000, 16} ;
}
